////////////////////////////////////////////////////////////////////////////////////////////////////

`include "encoder.vh"

////////////////////////////////////////////////////////////////////////////////////////////////////

module enc_par_buffer (
    input clk,
    input rst_n,
    input pro_finish,
    input [RSC_PAR_LEN - 1 : 0][EGF_DIM - 1 : 0] pro_data,
    output logic [ENC_PAR_BUF_DEP - 1 : 0][EGF_DIM - 1 : 0] par_buf_data
);

////////////////////////////////////////////////////////////////////////////////////////////////////

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            par_buf_data <= '0;
        end else if (pro_finish) begin
            par_buf_data <= pro_data;
        end
    end

endmodule

////////////////////////////////////////////////////////////////////////////////////////////////////