////////////////////////////////////////////////////////////////////////////////////////////////////

`include "encoder.vh"

////////////////////////////////////////////////////////////////////////////////////////////////////

module enc_mes_buffer (
    input clk,
    input rst_n,
    input con_stall,
    input [ENC_SYM - 1 : 0][EGF_DIM - 1 : 0] gen_data,
    output logic [ENC_MES_BUF_DEP - 1 : 0][EGF_DIM - 1 : 0] mes_buf_data
);

////////////////////////////////////////////////////////////////////////////////////////////////////

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            mes_buf_data <= '0;
        end else if (!con_stall) begin
            mes_buf_data[ENC_SYM - 1 : 0] <= gen_data;
            mes_buf_data[ENC_MES_BUF_DEP - 1 : ENC_SYM] <= mes_buf_data[ENC_MES_BUF_DEP - ENC_SYM - 1: 0];
        end
    end

endmodule

////////////////////////////////////////////////////////////////////////////////////////////////////